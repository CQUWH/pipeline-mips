// CQUWH
// 2020-12-25
`include "defines.vh"

module if_stage (
    
);

endmodule //if_stage