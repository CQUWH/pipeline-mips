// CQUWH
// 2020-12-25

module id_ex (
    
);

endmodule //id_ex