// CQUWH
// 2020-12-25
`include "defines.vh"

module mem_wb (
    
);

endmodule //mem_wb