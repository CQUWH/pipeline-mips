// CQUWH
// 2020-12-25

module main_decoder (
    
);

endmodule //main_decoder