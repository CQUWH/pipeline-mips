// CQUWH
// 2020-12-25

module ex_mem (
    
);

endmodule //ex_mem