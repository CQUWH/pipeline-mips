// CQUWH
// 2020-12-25

module branch_decoder (
    
);

endmodule //branch_decoder